library ieee; 

	-- STD_LOGIC and STD_LOGIC_VECTOR types, and relevant functions
	use ieee.std_logic_1164.all;

	-- SIGNED and UNSIGNED types, and relevant functions
	use ieee.numeric_std.all;
entity proyect2 is
	port (
		input : in std_LOGIC
	);
end entity;

architecture arch of proyect2 is

begin

end architecture;